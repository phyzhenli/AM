`timescale 1ns/1ps

module optimal3(
    input  [7:0]  x,
    input  [7:0]  y,
    output [15:0] z
);

wire [15:0] x0 = x << 7;
wire [15:0] y0 = y << 7;
wire signed [16:0] z0 = $signed(x0) + $signed(y0) - 16384;

wire [16:0] x_wire = x;
wire [16:0] y_wire = y;

wire signed [16:0] detz1 = (x>=0 && x<128 && y>=0 && y<128)? ($signed(x_wire))*(64-128)+($signed(y_wire))*(64-128)+128*128-64*64
: (x>=0 && x<128 && y>=128 && y<256)? ($signed(x_wire))*(192-128)+($signed(y_wire))*(64-128)+128*128-64*192
: (x>=128 && x<256 && y>=0 && y<128)? ($signed(x_wire))*(64-128)+($signed(y_wire))*(192-128)+128*128-192*64
: (x>=128 && x<256 && y>=128 && y<256)? ($signed(x_wire))*(192-128)+($signed(y_wire))*(192-128)+128*128-192*192
: 0;

wire signed [16:0] detz2 = (x>=0 && x<64 && y>=0 && y<64)? ($signed(x_wire))*(32-64)+($signed(y_wire))*(32-64)+64*64-32*32
: (x>=0 && x<64 && y>=64 && y<128)? ($signed(x_wire))*(96-64)+($signed(y_wire))*(32-64)+64*64-32*96
: (x>=0 && x<64 && y>=128 && y<192)? ($signed(x_wire))*(160-192)+($signed(y_wire))*(32-64)+64*192-32*160
: (x>=0 && x<64 && y>=192 && y<256)? ($signed(x_wire))*(224-192)+($signed(y_wire))*(32-64)+64*192-32*224
: (x>=64 && x<128 && y>=0 && y<64)? ($signed(x_wire))*(32-64)+($signed(y_wire))*(96-64)+64*64-96*32
: (x>=64 && x<128 && y>=64 && y<128)? ($signed(x_wire))*(96-64)+($signed(y_wire))*(96-64)+64*64-96*96
: (x>=64 && x<128 && y>=128 && y<192)? ($signed(x_wire))*(160-192)+($signed(y_wire))*(96-64)+64*192-96*160
: (x>=64 && x<128 && y>=192 && y<256)? ($signed(x_wire))*(224-192)+($signed(y_wire))*(96-64)+64*192-96*224
: (x>=128 && x<192 && y>=0 && y<64)? ($signed(x_wire))*(32-64)+($signed(y_wire))*(160-192)+192*64-160*32
: (x>=128 && x<192 && y>=64 && y<128)? ($signed(x_wire))*(96-64)+($signed(y_wire))*(160-192)+192*64-160*96
: (x>=128 && x<192 && y>=128 && y<192)? ($signed(x_wire))*(160-192)+($signed(y_wire))*(160-192)+192*192-160*160
: (x>=128 && x<192 && y>=192 && y<256)? ($signed(x_wire))*(224-192)+($signed(y_wire))*(160-192)+192*192-160*224
: (x>=192 && x<256 && y>=0 && y<64)? ($signed(x_wire))*(32-64)+($signed(y_wire))*(224-192)+192*64-224*32
: (x>=192 && x<256 && y>=64 && y<128)? ($signed(x_wire))*(96-64)+($signed(y_wire))*(224-192)+192*64-224*96
: (x>=192 && x<256 && y>=128 && y<192)? ($signed(x_wire))*(160-192)+($signed(y_wire))*(224-192)+192*192-224*160
: (x>=192 && x<256 && y>=192 && y<256)? ($signed(x_wire))*(224-192)+($signed(y_wire))*(224-192)+192*192-224*224
: 0;


wire signed [16:0] detz3 = (x>=0 && x<32 && y>=0 && y<32)? ($signed(x_wire))*(16-32)+($signed(y_wire))*(16-32)+32*32-16*16
: (x>=0 && x<32 && y>=32 && y<64)? ($signed(x_wire))*(48-32)+($signed(y_wire))*(16-32)+32*32-16*48
: (x>=0 && x<32 && y>=64 && y<96)? ($signed(x_wire))*(80-96)+($signed(y_wire))*(16-32)+32*96-16*80
: (x>=0 && x<32 && y>=96 && y<128)? ($signed(x_wire))*(112-96)+($signed(y_wire))*(16-32)+32*96-16*112
: (x>=0 && x<32 && y>=128 && y<160)? ($signed(x_wire))*(144-160)+($signed(y_wire))*(16-32)+32*160-16*144
: (x>=0 && x<32 && y>=160 && y<192)? ($signed(x_wire))*(176-160)+($signed(y_wire))*(16-32)+32*160-16*176
: (x>=0 && x<32 && y>=192 && y<224)? ($signed(x_wire))*(208-224)+($signed(y_wire))*(16-32)+32*224-16*208
: (x>=0 && x<32 && y>=224 && y<256)? ($signed(x_wire))*(240-224)+($signed(y_wire))*(16-32)+32*224-16*240
: (x>=32 && x<64 && y>=0 && y<32)? ($signed(x_wire))*(16-32)+($signed(y_wire))*(48-32)+32*32-48*16
: (x>=32 && x<64 && y>=32 && y<64)? ($signed(x_wire))*(48-32)+($signed(y_wire))*(48-32)+32*32-48*48
: (x>=32 && x<64 && y>=64 && y<96)? ($signed(x_wire))*(80-96)+($signed(y_wire))*(48-32)+32*96-48*80
: (x>=32 && x<64 && y>=96 && y<128)? ($signed(x_wire))*(112-96)+($signed(y_wire))*(48-32)+32*96-48*112
: (x>=32 && x<64 && y>=128 && y<160)? ($signed(x_wire))*(144-160)+($signed(y_wire))*(48-32)+32*160-48*144
: (x>=32 && x<64 && y>=160 && y<192)? ($signed(x_wire))*(176-160)+($signed(y_wire))*(48-32)+32*160-48*176
: (x>=32 && x<64 && y>=192 && y<224)? ($signed(x_wire))*(208-224)+($signed(y_wire))*(48-32)+32*224-48*208
: (x>=32 && x<64 && y>=224 && y<256)? ($signed(x_wire))*(240-224)+($signed(y_wire))*(48-32)+32*224-48*240
: (x>=64 && x<96 && y>=0 && y<32)? ($signed(x_wire))*(16-32)+($signed(y_wire))*(80-96)+96*32-80*16
: (x>=64 && x<96 && y>=32 && y<64)? ($signed(x_wire))*(48-32)+($signed(y_wire))*(80-96)+96*32-80*48
: (x>=64 && x<96 && y>=64 && y<96)? ($signed(x_wire))*(80-96)+($signed(y_wire))*(80-96)+96*96-80*80
: (x>=64 && x<96 && y>=96 && y<128)? ($signed(x_wire))*(112-96)+($signed(y_wire))*(80-96)+96*96-80*112
: (x>=64 && x<96 && y>=128 && y<160)? ($signed(x_wire))*(144-160)+($signed(y_wire))*(80-96)+96*160-80*144
: (x>=64 && x<96 && y>=160 && y<192)? ($signed(x_wire))*(176-160)+($signed(y_wire))*(80-96)+96*160-80*176
: (x>=64 && x<96 && y>=192 && y<224)? ($signed(x_wire))*(208-224)+($signed(y_wire))*(80-96)+96*224-80*208
: (x>=64 && x<96 && y>=224 && y<256)? ($signed(x_wire))*(240-224)+($signed(y_wire))*(80-96)+96*224-80*240
: (x>=96 && x<128 && y>=0 && y<32)? ($signed(x_wire))*(16-32)+($signed(y_wire))*(112-96)+96*32-112*16
: (x>=96 && x<128 && y>=32 && y<64)? ($signed(x_wire))*(48-32)+($signed(y_wire))*(112-96)+96*32-112*48
: (x>=96 && x<128 && y>=64 && y<96)? ($signed(x_wire))*(80-96)+($signed(y_wire))*(112-96)+96*96-112*80
: (x>=96 && x<128 && y>=96 && y<128)? ($signed(x_wire))*(112-96)+($signed(y_wire))*(112-96)+96*96-112*112
: (x>=96 && x<128 && y>=128 && y<160)? ($signed(x_wire))*(144-160)+($signed(y_wire))*(112-96)+96*160-112*144
: (x>=96 && x<128 && y>=160 && y<192)? ($signed(x_wire))*(176-160)+($signed(y_wire))*(112-96)+96*160-112*176
: (x>=96 && x<128 && y>=192 && y<224)? ($signed(x_wire))*(208-224)+($signed(y_wire))*(112-96)+96*224-112*208
: (x>=96 && x<128 && y>=224 && y<256)? ($signed(x_wire))*(240-224)+($signed(y_wire))*(112-96)+96*224-112*240
: (x>=128 && x<160 && y>=0 && y<32)? ($signed(x_wire))*(16-32)+($signed(y_wire))*(144-160)+160*32-144*16
: (x>=128 && x<160 && y>=32 && y<64)? ($signed(x_wire))*(48-32)+($signed(y_wire))*(144-160)+160*32-144*48
: (x>=128 && x<160 && y>=64 && y<96)? ($signed(x_wire))*(80-96)+($signed(y_wire))*(144-160)+160*96-144*80
: (x>=128 && x<160 && y>=96 && y<128)? ($signed(x_wire))*(112-96)+($signed(y_wire))*(144-160)+160*96-144*112
: (x>=128 && x<160 && y>=128 && y<160)? ($signed(x_wire))*(144-160)+($signed(y_wire))*(144-160)+160*160-144*144
: (x>=128 && x<160 && y>=160 && y<192)? ($signed(x_wire))*(176-160)+($signed(y_wire))*(144-160)+160*160-144*176
: (x>=128 && x<160 && y>=192 && y<224)? ($signed(x_wire))*(208-224)+($signed(y_wire))*(144-160)+160*224-144*208
: (x>=128 && x<160 && y>=224 && y<256)? ($signed(x_wire))*(240-224)+($signed(y_wire))*(144-160)+160*224-144*240
: (x>=160 && x<192 && y>=0 && y<32)? ($signed(x_wire))*(16-32)+($signed(y_wire))*(176-160)+160*32-176*16
: (x>=160 && x<192 && y>=32 && y<64)? ($signed(x_wire))*(48-32)+($signed(y_wire))*(176-160)+160*32-176*48
: (x>=160 && x<192 && y>=64 && y<96)? ($signed(x_wire))*(80-96)+($signed(y_wire))*(176-160)+160*96-176*80
: (x>=160 && x<192 && y>=96 && y<128)? ($signed(x_wire))*(112-96)+($signed(y_wire))*(176-160)+160*96-176*112
: (x>=160 && x<192 && y>=128 && y<160)? ($signed(x_wire))*(144-160)+($signed(y_wire))*(176-160)+160*160-176*144
: (x>=160 && x<192 && y>=160 && y<192)? ($signed(x_wire))*(176-160)+($signed(y_wire))*(176-160)+160*160-176*176
: (x>=160 && x<192 && y>=192 && y<224)? ($signed(x_wire))*(208-224)+($signed(y_wire))*(176-160)+160*224-176*208
: (x>=160 && x<192 && y>=224 && y<256)? ($signed(x_wire))*(240-224)+($signed(y_wire))*(176-160)+160*224-176*240
: (x>=192 && x<224 && y>=0 && y<32)? ($signed(x_wire))*(16-32)+($signed(y_wire))*(208-224)+224*32-208*16
: (x>=192 && x<224 && y>=32 && y<64)? ($signed(x_wire))*(48-32)+($signed(y_wire))*(208-224)+224*32-208*48
: (x>=192 && x<224 && y>=64 && y<96)? ($signed(x_wire))*(80-96)+($signed(y_wire))*(208-224)+224*96-208*80
: (x>=192 && x<224 && y>=96 && y<128)? ($signed(x_wire))*(112-96)+($signed(y_wire))*(208-224)+224*96-208*112
: (x>=192 && x<224 && y>=128 && y<160)? ($signed(x_wire))*(144-160)+($signed(y_wire))*(208-224)+224*160-208*144
: (x>=192 && x<224 && y>=160 && y<192)? ($signed(x_wire))*(176-160)+($signed(y_wire))*(208-224)+224*160-208*176
: (x>=192 && x<224 && y>=192 && y<224)? ($signed(x_wire))*(208-224)+($signed(y_wire))*(208-224)+224*224-208*208
: (x>=192 && x<224 && y>=224 && y<256)? ($signed(x_wire))*(240-224)+($signed(y_wire))*(208-224)+224*224-208*240
: (x>=224 && x<256 && y>=0 && y<32)? ($signed(x_wire))*(16-32)+($signed(y_wire))*(240-224)+224*32-240*16
: (x>=224 && x<256 && y>=32 && y<64)? ($signed(x_wire))*(48-32)+($signed(y_wire))*(240-224)+224*32-240*48
: (x>=224 && x<256 && y>=64 && y<96)? ($signed(x_wire))*(80-96)+($signed(y_wire))*(240-224)+224*96-240*80
: (x>=224 && x<256 && y>=96 && y<128)? ($signed(x_wire))*(112-96)+($signed(y_wire))*(240-224)+224*96-240*112
: (x>=224 && x<256 && y>=128 && y<160)? ($signed(x_wire))*(144-160)+($signed(y_wire))*(240-224)+224*160-240*144
: (x>=224 && x<256 && y>=160 && y<192)? ($signed(x_wire))*(176-160)+($signed(y_wire))*(240-224)+224*160-240*176
: (x>=224 && x<256 && y>=192 && y<224)? ($signed(x_wire))*(208-224)+($signed(y_wire))*(240-224)+224*224-240*208
: (x>=224 && x<256 && y>=224 && y<256)? ($signed(x_wire))*(240-224)+($signed(y_wire))*(240-224)+224*224-240*240
: 0;

wire signed [16:0] detz4 = (x>=0 && x<16 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(8-16)+16*16-8*8
: (x>=0 && x<16 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(8-16)+16*16-8*24
: (x>=0 && x<16 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(8-16)+16*48-8*40
: (x>=0 && x<16 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(8-16)+16*48-8*56
: (x>=0 && x<16 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(8-16)+16*80-8*72
: (x>=0 && x<16 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(8-16)+16*80-8*88
: (x>=0 && x<16 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(8-16)+16*112-8*104
: (x>=0 && x<16 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(8-16)+16*112-8*120
: (x>=0 && x<16 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(8-16)+16*144-8*136
: (x>=0 && x<16 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(8-16)+16*144-8*152
: (x>=0 && x<16 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(8-16)+16*176-8*168
: (x>=0 && x<16 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(8-16)+16*176-8*184
: (x>=0 && x<16 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(8-16)+16*208-8*200
: (x>=0 && x<16 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(8-16)+16*208-8*216
: (x>=0 && x<16 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(8-16)+16*240-8*232
: (x>=0 && x<16 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(8-16)+16*240-8*248
: (x>=16 && x<32 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(24-16)+16*16-24*8
: (x>=16 && x<32 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(24-16)+16*16-24*24
: (x>=16 && x<32 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(24-16)+16*48-24*40
: (x>=16 && x<32 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(24-16)+16*48-24*56
: (x>=16 && x<32 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(24-16)+16*80-24*72
: (x>=16 && x<32 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(24-16)+16*80-24*88
: (x>=16 && x<32 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(24-16)+16*112-24*104
: (x>=16 && x<32 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(24-16)+16*112-24*120
: (x>=16 && x<32 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(24-16)+16*144-24*136
: (x>=16 && x<32 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(24-16)+16*144-24*152
: (x>=16 && x<32 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(24-16)+16*176-24*168
: (x>=16 && x<32 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(24-16)+16*176-24*184
: (x>=16 && x<32 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(24-16)+16*208-24*200
: (x>=16 && x<32 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(24-16)+16*208-24*216
: (x>=16 && x<32 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(24-16)+16*240-24*232
: (x>=16 && x<32 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(24-16)+16*240-24*248
: (x>=32 && x<48 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(40-48)+48*16-40*8
: (x>=32 && x<48 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(40-48)+48*16-40*24
: (x>=32 && x<48 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(40-48)+48*48-40*40
: (x>=32 && x<48 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(40-48)+48*48-40*56
: (x>=32 && x<48 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(40-48)+48*80-40*72
: (x>=32 && x<48 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(40-48)+48*80-40*88
: (x>=32 && x<48 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(40-48)+48*112-40*104
: (x>=32 && x<48 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(40-48)+48*112-40*120
: (x>=32 && x<48 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(40-48)+48*144-40*136
: (x>=32 && x<48 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(40-48)+48*144-40*152
: (x>=32 && x<48 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(40-48)+48*176-40*168
: (x>=32 && x<48 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(40-48)+48*176-40*184
: (x>=32 && x<48 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(40-48)+48*208-40*200
: (x>=32 && x<48 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(40-48)+48*208-40*216
: (x>=32 && x<48 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(40-48)+48*240-40*232
: (x>=32 && x<48 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(40-48)+48*240-40*248
: (x>=48 && x<64 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(56-48)+48*16-56*8
: (x>=48 && x<64 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(56-48)+48*16-56*24
: (x>=48 && x<64 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(56-48)+48*48-56*40
: (x>=48 && x<64 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(56-48)+48*48-56*56
: (x>=48 && x<64 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(56-48)+48*80-56*72
: (x>=48 && x<64 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(56-48)+48*80-56*88
: (x>=48 && x<64 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(56-48)+48*112-56*104
: (x>=48 && x<64 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(56-48)+48*112-56*120
: (x>=48 && x<64 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(56-48)+48*144-56*136
: (x>=48 && x<64 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(56-48)+48*144-56*152
: (x>=48 && x<64 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(56-48)+48*176-56*168
: (x>=48 && x<64 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(56-48)+48*176-56*184
: (x>=48 && x<64 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(56-48)+48*208-56*200
: (x>=48 && x<64 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(56-48)+48*208-56*216
: (x>=48 && x<64 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(56-48)+48*240-56*232
: (x>=48 && x<64 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(56-48)+48*240-56*248
: (x>=64 && x<80 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(72-80)+80*16-72*8
: (x>=64 && x<80 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(72-80)+80*16-72*24
: (x>=64 && x<80 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(72-80)+80*48-72*40
: (x>=64 && x<80 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(72-80)+80*48-72*56
: (x>=64 && x<80 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(72-80)+80*80-72*72
: (x>=64 && x<80 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(72-80)+80*80-72*88
: (x>=64 && x<80 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(72-80)+80*112-72*104
: (x>=64 && x<80 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(72-80)+80*112-72*120
: (x>=64 && x<80 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(72-80)+80*144-72*136
: (x>=64 && x<80 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(72-80)+80*144-72*152
: (x>=64 && x<80 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(72-80)+80*176-72*168
: (x>=64 && x<80 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(72-80)+80*176-72*184
: (x>=64 && x<80 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(72-80)+80*208-72*200
: (x>=64 && x<80 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(72-80)+80*208-72*216
: (x>=64 && x<80 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(72-80)+80*240-72*232
: (x>=64 && x<80 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(72-80)+80*240-72*248
: (x>=80 && x<96 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(88-80)+80*16-88*8
: (x>=80 && x<96 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(88-80)+80*16-88*24
: (x>=80 && x<96 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(88-80)+80*48-88*40
: (x>=80 && x<96 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(88-80)+80*48-88*56
: (x>=80 && x<96 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(88-80)+80*80-88*72
: (x>=80 && x<96 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(88-80)+80*80-88*88
: (x>=80 && x<96 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(88-80)+80*112-88*104
: (x>=80 && x<96 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(88-80)+80*112-88*120
: (x>=80 && x<96 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(88-80)+80*144-88*136
: (x>=80 && x<96 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(88-80)+80*144-88*152
: (x>=80 && x<96 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(88-80)+80*176-88*168
: (x>=80 && x<96 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(88-80)+80*176-88*184
: (x>=80 && x<96 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(88-80)+80*208-88*200
: (x>=80 && x<96 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(88-80)+80*208-88*216
: (x>=80 && x<96 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(88-80)+80*240-88*232
: (x>=80 && x<96 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(88-80)+80*240-88*248
: (x>=96 && x<112 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(104-112)+112*16-104*8
: (x>=96 && x<112 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(104-112)+112*16-104*24
: (x>=96 && x<112 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(104-112)+112*48-104*40
: (x>=96 && x<112 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(104-112)+112*48-104*56
: (x>=96 && x<112 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(104-112)+112*80-104*72
: (x>=96 && x<112 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(104-112)+112*80-104*88
: (x>=96 && x<112 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(104-112)+112*112-104*104
: (x>=96 && x<112 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(104-112)+112*112-104*120
: (x>=96 && x<112 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(104-112)+112*144-104*136
: (x>=96 && x<112 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(104-112)+112*144-104*152
: (x>=96 && x<112 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(104-112)+112*176-104*168
: (x>=96 && x<112 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(104-112)+112*176-104*184
: (x>=96 && x<112 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(104-112)+112*208-104*200
: (x>=96 && x<112 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(104-112)+112*208-104*216
: (x>=96 && x<112 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(104-112)+112*240-104*232
: (x>=96 && x<112 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(104-112)+112*240-104*248
: (x>=112 && x<128 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(120-112)+112*16-120*8
: (x>=112 && x<128 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(120-112)+112*16-120*24
: (x>=112 && x<128 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(120-112)+112*48-120*40
: (x>=112 && x<128 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(120-112)+112*48-120*56
: (x>=112 && x<128 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(120-112)+112*80-120*72
: (x>=112 && x<128 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(120-112)+112*80-120*88
: (x>=112 && x<128 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(120-112)+112*112-120*104
: (x>=112 && x<128 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(120-112)+112*112-120*120
: (x>=112 && x<128 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(120-112)+112*144-120*136
: (x>=112 && x<128 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(120-112)+112*144-120*152
: (x>=112 && x<128 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(120-112)+112*176-120*168
: (x>=112 && x<128 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(120-112)+112*176-120*184
: (x>=112 && x<128 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(120-112)+112*208-120*200
: (x>=112 && x<128 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(120-112)+112*208-120*216
: (x>=112 && x<128 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(120-112)+112*240-120*232
: (x>=112 && x<128 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(120-112)+112*240-120*248
: (x>=128 && x<144 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(136-144)+144*16-136*8
: (x>=128 && x<144 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(136-144)+144*16-136*24
: (x>=128 && x<144 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(136-144)+144*48-136*40
: (x>=128 && x<144 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(136-144)+144*48-136*56
: (x>=128 && x<144 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(136-144)+144*80-136*72
: (x>=128 && x<144 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(136-144)+144*80-136*88
: (x>=128 && x<144 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(136-144)+144*112-136*104
: (x>=128 && x<144 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(136-144)+144*112-136*120
: (x>=128 && x<144 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(136-144)+144*144-136*136
: (x>=128 && x<144 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(136-144)+144*144-136*152
: (x>=128 && x<144 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(136-144)+144*176-136*168
: (x>=128 && x<144 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(136-144)+144*176-136*184
: (x>=128 && x<144 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(136-144)+144*208-136*200
: (x>=128 && x<144 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(136-144)+144*208-136*216
: (x>=128 && x<144 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(136-144)+144*240-136*232
: (x>=128 && x<144 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(136-144)+144*240-136*248
: (x>=144 && x<160 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(152-144)+144*16-152*8
: (x>=144 && x<160 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(152-144)+144*16-152*24
: (x>=144 && x<160 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(152-144)+144*48-152*40
: (x>=144 && x<160 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(152-144)+144*48-152*56
: (x>=144 && x<160 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(152-144)+144*80-152*72
: (x>=144 && x<160 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(152-144)+144*80-152*88
: (x>=144 && x<160 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(152-144)+144*112-152*104
: (x>=144 && x<160 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(152-144)+144*112-152*120
: (x>=144 && x<160 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(152-144)+144*144-152*136
: (x>=144 && x<160 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(152-144)+144*144-152*152
: (x>=144 && x<160 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(152-144)+144*176-152*168
: (x>=144 && x<160 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(152-144)+144*176-152*184
: (x>=144 && x<160 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(152-144)+144*208-152*200
: (x>=144 && x<160 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(152-144)+144*208-152*216
: (x>=144 && x<160 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(152-144)+144*240-152*232
: (x>=144 && x<160 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(152-144)+144*240-152*248
: (x>=160 && x<176 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(168-176)+176*16-168*8
: (x>=160 && x<176 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(168-176)+176*16-168*24
: (x>=160 && x<176 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(168-176)+176*48-168*40
: (x>=160 && x<176 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(168-176)+176*48-168*56
: (x>=160 && x<176 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(168-176)+176*80-168*72
: (x>=160 && x<176 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(168-176)+176*80-168*88
: (x>=160 && x<176 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(168-176)+176*112-168*104
: (x>=160 && x<176 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(168-176)+176*112-168*120
: (x>=160 && x<176 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(168-176)+176*144-168*136
: (x>=160 && x<176 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(168-176)+176*144-168*152
: (x>=160 && x<176 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(168-176)+176*176-168*168
: (x>=160 && x<176 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(168-176)+176*176-168*184
: (x>=160 && x<176 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(168-176)+176*208-168*200
: (x>=160 && x<176 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(168-176)+176*208-168*216
: (x>=160 && x<176 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(168-176)+176*240-168*232
: (x>=160 && x<176 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(168-176)+176*240-168*248
: (x>=176 && x<192 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(184-176)+176*16-184*8
: (x>=176 && x<192 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(184-176)+176*16-184*24
: (x>=176 && x<192 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(184-176)+176*48-184*40
: (x>=176 && x<192 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(184-176)+176*48-184*56
: (x>=176 && x<192 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(184-176)+176*80-184*72
: (x>=176 && x<192 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(184-176)+176*80-184*88
: (x>=176 && x<192 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(184-176)+176*112-184*104
: (x>=176 && x<192 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(184-176)+176*112-184*120
: (x>=176 && x<192 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(184-176)+176*144-184*136
: (x>=176 && x<192 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(184-176)+176*144-184*152
: (x>=176 && x<192 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(184-176)+176*176-184*168
: (x>=176 && x<192 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(184-176)+176*176-184*184
: (x>=176 && x<192 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(184-176)+176*208-184*200
: (x>=176 && x<192 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(184-176)+176*208-184*216
: (x>=176 && x<192 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(184-176)+176*240-184*232
: (x>=176 && x<192 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(184-176)+176*240-184*248
: (x>=192 && x<208 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(200-208)+208*16-200*8
: (x>=192 && x<208 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(200-208)+208*16-200*24
: (x>=192 && x<208 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(200-208)+208*48-200*40
: (x>=192 && x<208 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(200-208)+208*48-200*56
: (x>=192 && x<208 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(200-208)+208*80-200*72
: (x>=192 && x<208 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(200-208)+208*80-200*88
: (x>=192 && x<208 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(200-208)+208*112-200*104
: (x>=192 && x<208 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(200-208)+208*112-200*120
: (x>=192 && x<208 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(200-208)+208*144-200*136
: (x>=192 && x<208 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(200-208)+208*144-200*152
: (x>=192 && x<208 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(200-208)+208*176-200*168
: (x>=192 && x<208 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(200-208)+208*176-200*184
: (x>=192 && x<208 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(200-208)+208*208-200*200
: (x>=192 && x<208 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(200-208)+208*208-200*216
: (x>=192 && x<208 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(200-208)+208*240-200*232
: (x>=192 && x<208 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(200-208)+208*240-200*248
: (x>=208 && x<224 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(216-208)+208*16-216*8
: (x>=208 && x<224 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(216-208)+208*16-216*24
: (x>=208 && x<224 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(216-208)+208*48-216*40
: (x>=208 && x<224 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(216-208)+208*48-216*56
: (x>=208 && x<224 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(216-208)+208*80-216*72
: (x>=208 && x<224 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(216-208)+208*80-216*88
: (x>=208 && x<224 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(216-208)+208*112-216*104
: (x>=208 && x<224 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(216-208)+208*112-216*120
: (x>=208 && x<224 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(216-208)+208*144-216*136
: (x>=208 && x<224 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(216-208)+208*144-216*152
: (x>=208 && x<224 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(216-208)+208*176-216*168
: (x>=208 && x<224 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(216-208)+208*176-216*184
: (x>=208 && x<224 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(216-208)+208*208-216*200
: (x>=208 && x<224 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(216-208)+208*208-216*216
: (x>=208 && x<224 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(216-208)+208*240-216*232
: (x>=208 && x<224 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(216-208)+208*240-216*248
: (x>=224 && x<240 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(232-240)+240*16-232*8
: (x>=224 && x<240 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(232-240)+240*16-232*24
: (x>=224 && x<240 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(232-240)+240*48-232*40
: (x>=224 && x<240 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(232-240)+240*48-232*56
: (x>=224 && x<240 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(232-240)+240*80-232*72
: (x>=224 && x<240 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(232-240)+240*80-232*88
: (x>=224 && x<240 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(232-240)+240*112-232*104
: (x>=224 && x<240 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(232-240)+240*112-232*120
: (x>=224 && x<240 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(232-240)+240*144-232*136
: (x>=224 && x<240 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(232-240)+240*144-232*152
: (x>=224 && x<240 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(232-240)+240*176-232*168
: (x>=224 && x<240 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(232-240)+240*176-232*184
: (x>=224 && x<240 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(232-240)+240*208-232*200
: (x>=224 && x<240 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(232-240)+240*208-232*216
: (x>=224 && x<240 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(232-240)+240*240-232*232
: (x>=224 && x<240 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(232-240)+240*240-232*248
: (x>=240 && x<256 && y>=0 && y<16)? ($signed(x_wire))*(8-16)+($signed(y_wire))*(248-240)+240*16-248*8
: (x>=240 && x<256 && y>=16 && y<32)? ($signed(x_wire))*(24-16)+($signed(y_wire))*(248-240)+240*16-248*24
: (x>=240 && x<256 && y>=32 && y<48)? ($signed(x_wire))*(40-48)+($signed(y_wire))*(248-240)+240*48-248*40
: (x>=240 && x<256 && y>=48 && y<64)? ($signed(x_wire))*(56-48)+($signed(y_wire))*(248-240)+240*48-248*56
: (x>=240 && x<256 && y>=64 && y<80)? ($signed(x_wire))*(72-80)+($signed(y_wire))*(248-240)+240*80-248*72
: (x>=240 && x<256 && y>=80 && y<96)? ($signed(x_wire))*(88-80)+($signed(y_wire))*(248-240)+240*80-248*88
: (x>=240 && x<256 && y>=96 && y<112)? ($signed(x_wire))*(104-112)+($signed(y_wire))*(248-240)+240*112-248*104
: (x>=240 && x<256 && y>=112 && y<128)? ($signed(x_wire))*(120-112)+($signed(y_wire))*(248-240)+240*112-248*120
: (x>=240 && x<256 && y>=128 && y<144)? ($signed(x_wire))*(136-144)+($signed(y_wire))*(248-240)+240*144-248*136
: (x>=240 && x<256 && y>=144 && y<160)? ($signed(x_wire))*(152-144)+($signed(y_wire))*(248-240)+240*144-248*152
: (x>=240 && x<256 && y>=160 && y<176)? ($signed(x_wire))*(168-176)+($signed(y_wire))*(248-240)+240*176-248*168
: (x>=240 && x<256 && y>=176 && y<192)? ($signed(x_wire))*(184-176)+($signed(y_wire))*(248-240)+240*176-248*184
: (x>=240 && x<256 && y>=192 && y<208)? ($signed(x_wire))*(200-208)+($signed(y_wire))*(248-240)+240*208-248*200
: (x>=240 && x<256 && y>=208 && y<224)? ($signed(x_wire))*(216-208)+($signed(y_wire))*(248-240)+240*208-248*216
: (x>=240 && x<256 && y>=224 && y<240)? ($signed(x_wire))*(232-240)+($signed(y_wire))*(248-240)+240*240-248*232
: (x>=240 && x<256 && y>=240 && y<256)? ($signed(x_wire))*(248-240)+($signed(y_wire))*(248-240)+240*240-248*248
: 0;

wire signed [16:0] z_sign = z0 + detz1 + detz2 + detz3;

assign z = (z_sign < 0)? 0 : z_sign[15:0];

endmodule
