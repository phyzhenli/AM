module ubit8_designware(input [7:0] a1,b1, output [15:0] result
    );
	 
	assign result = a1*b1;

endmodule
