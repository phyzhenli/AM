module FIFO(
  input        clock,
  input        reset,
  input  [7:0] io_din,
  input        io_wr_en,
  input        io_rd_en,
  output       io_empty,
  output [7:0] io_dout
);
  reg [7:0] mem_0; // @[fifo.scala 15:22]
  reg [31:0] _RAND_0;
  reg [7:0] mem_1; // @[fifo.scala 15:22]
  reg [31:0] _RAND_1;
  reg [7:0] mem_2; // @[fifo.scala 15:22]
  reg [31:0] _RAND_2;
  reg [7:0] mem_3; // @[fifo.scala 15:22]
  reg [31:0] _RAND_3;
  reg [7:0] mem_4; // @[fifo.scala 15:22]
  reg [31:0] _RAND_4;
  reg [7:0] mem_5; // @[fifo.scala 15:22]
  reg [31:0] _RAND_5;
  reg [7:0] mem_6; // @[fifo.scala 15:22]
  reg [31:0] _RAND_6;
  reg [7:0] mem_7; // @[fifo.scala 15:22]
  reg [31:0] _RAND_7;
  reg [7:0] mem_8; // @[fifo.scala 15:22]
  reg [31:0] _RAND_8;
  reg [7:0] mem_9; // @[fifo.scala 15:22]
  reg [31:0] _RAND_9;
  reg [7:0] mem_10; // @[fifo.scala 15:22]
  reg [31:0] _RAND_10;
  reg [7:0] mem_11; // @[fifo.scala 15:22]
  reg [31:0] _RAND_11;
  reg [7:0] mem_12; // @[fifo.scala 15:22]
  reg [31:0] _RAND_12;
  reg [7:0] mem_13; // @[fifo.scala 15:22]
  reg [31:0] _RAND_13;
  reg [7:0] mem_14; // @[fifo.scala 15:22]
  reg [31:0] _RAND_14;
  reg [7:0] mem_15; // @[fifo.scala 15:22]
  reg [31:0] _RAND_15;
  reg [7:0] dout_reg; // @[fifo.scala 17:27]
  reg [31:0] _RAND_16;
  reg  empty_reg; // @[fifo.scala 18:28]
  reg [31:0] _RAND_17;
  reg [3:0] wr_sp; // @[fifo.scala 22:24]
  reg [31:0] _RAND_18;
  wire  _T_1; // @[fifo.scala 25:22]
  wire  _T_2; // @[fifo.scala 25:19]
  wire [3:0] _T_4; // @[fifo.scala 26:24]
  wire  _GEN_33; // @[fifo.scala 25:33]
  wire  _T_5; // @[fifo.scala 31:10]
  wire  _T_6; // @[fifo.scala 31:20]
  wire  _T_7; // @[fifo.scala 32:20]
  wire [3:0] _T_9; // @[fifo.scala 34:28]
  wire  _T_10; // @[fifo.scala 41:25]
  wire  _GEN_68; // @[fifo.scala 32:37]
  wire  _GEN_87; // @[fifo.scala 31:33]
  wire  _T_13; // @[fifo.scala 52:19]
  wire [4:0] _GEN_176; // @[fifo.scala 53:20]
  wire  _T_14; // @[fifo.scala 53:20]
  wire  _GEN_155; // @[fifo.scala 54:9]
  wire  _GEN_174; // @[fifo.scala 52:32]
  assign _T_1 = io_rd_en == 1'h0; // @[fifo.scala 25:22]
  assign _T_2 = io_wr_en & _T_1; // @[fifo.scala 25:19]
  assign _T_4 = wr_sp - 4'h1; // @[fifo.scala 26:24]
  assign _GEN_33 = _T_2 ? 1'h0 : empty_reg; // @[fifo.scala 25:33]
  assign _T_5 = io_wr_en == 1'h0; // @[fifo.scala 31:10]
  assign _T_6 = _T_5 & io_rd_en; // @[fifo.scala 31:20]
  assign _T_7 = wr_sp == 4'he; // @[fifo.scala 32:20]
  assign _T_9 = wr_sp + 4'h1; // @[fifo.scala 34:28]
  assign _T_10 = wr_sp == 4'hf; // @[fifo.scala 41:25]
  assign _GEN_68 = _T_7 | _GEN_33; // @[fifo.scala 32:37]
  assign _GEN_87 = _T_6 ? _GEN_68 : _GEN_33; // @[fifo.scala 31:33]
  assign _T_13 = io_wr_en & io_rd_en; // @[fifo.scala 52:19]
  assign _GEN_176 = {{1'd0}, wr_sp}; // @[fifo.scala 53:20]
  assign _T_14 = _GEN_176 == 5'h10; // @[fifo.scala 53:20]
  assign _GEN_155 = _T_14 ? 1'h0 : _GEN_87; // @[fifo.scala 54:9]
  assign _GEN_174 = _T_13 ? _GEN_155 : _GEN_87; // @[fifo.scala 52:32]
  assign io_empty = empty_reg; // @[fifo.scala 20:14]
  assign io_dout = dout_reg; // @[fifo.scala 19:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  dout_reg = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  empty_reg = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wr_sp = _RAND_18[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      mem_0 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h0 == wr_sp) begin
            mem_0 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_0 <= 8'h0;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h0 == wr_sp) begin
                      mem_0 <= io_din;
                    end
                  end
                end else begin
                  mem_0 <= 8'h0;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h0 == wr_sp) begin
                  mem_0 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_0 <= 8'h0;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_0 <= 8'h0;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h0 == wr_sp) begin
                  mem_0 <= io_din;
                end
              end
            end else begin
              mem_0 <= 8'h0;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h0 == wr_sp) begin
              mem_0 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_1 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h1 == wr_sp) begin
            mem_1 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_1 <= mem_0;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h1 == wr_sp) begin
                      mem_1 <= io_din;
                    end
                  end
                end else begin
                  mem_1 <= mem_0;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h1 == wr_sp) begin
                  mem_1 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_1 <= mem_0;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_1 <= mem_0;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h1 == wr_sp) begin
                  mem_1 <= io_din;
                end
              end
            end else begin
              mem_1 <= mem_0;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h1 == wr_sp) begin
              mem_1 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_2 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h2 == wr_sp) begin
            mem_2 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_2 <= mem_1;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h2 == wr_sp) begin
                      mem_2 <= io_din;
                    end
                  end
                end else begin
                  mem_2 <= mem_1;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h2 == wr_sp) begin
                  mem_2 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_2 <= mem_1;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_2 <= mem_1;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h2 == wr_sp) begin
                  mem_2 <= io_din;
                end
              end
            end else begin
              mem_2 <= mem_1;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h2 == wr_sp) begin
              mem_2 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_3 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h3 == wr_sp) begin
            mem_3 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_3 <= mem_2;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h3 == wr_sp) begin
                      mem_3 <= io_din;
                    end
                  end
                end else begin
                  mem_3 <= mem_2;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h3 == wr_sp) begin
                  mem_3 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_3 <= mem_2;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_3 <= mem_2;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h3 == wr_sp) begin
                  mem_3 <= io_din;
                end
              end
            end else begin
              mem_3 <= mem_2;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h3 == wr_sp) begin
              mem_3 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_4 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h4 == wr_sp) begin
            mem_4 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_4 <= mem_3;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h4 == wr_sp) begin
                      mem_4 <= io_din;
                    end
                  end
                end else begin
                  mem_4 <= mem_3;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h4 == wr_sp) begin
                  mem_4 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_4 <= mem_3;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_4 <= mem_3;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h4 == wr_sp) begin
                  mem_4 <= io_din;
                end
              end
            end else begin
              mem_4 <= mem_3;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h4 == wr_sp) begin
              mem_4 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_5 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h5 == wr_sp) begin
            mem_5 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_5 <= mem_4;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h5 == wr_sp) begin
                      mem_5 <= io_din;
                    end
                  end
                end else begin
                  mem_5 <= mem_4;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h5 == wr_sp) begin
                  mem_5 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_5 <= mem_4;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_5 <= mem_4;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h5 == wr_sp) begin
                  mem_5 <= io_din;
                end
              end
            end else begin
              mem_5 <= mem_4;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h5 == wr_sp) begin
              mem_5 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_6 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h6 == wr_sp) begin
            mem_6 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_6 <= mem_5;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h6 == wr_sp) begin
                      mem_6 <= io_din;
                    end
                  end
                end else begin
                  mem_6 <= mem_5;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h6 == wr_sp) begin
                  mem_6 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_6 <= mem_5;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_6 <= mem_5;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h6 == wr_sp) begin
                  mem_6 <= io_din;
                end
              end
            end else begin
              mem_6 <= mem_5;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h6 == wr_sp) begin
              mem_6 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_7 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h7 == wr_sp) begin
            mem_7 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_7 <= mem_6;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h7 == wr_sp) begin
                      mem_7 <= io_din;
                    end
                  end
                end else begin
                  mem_7 <= mem_6;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h7 == wr_sp) begin
                  mem_7 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_7 <= mem_6;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_7 <= mem_6;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h7 == wr_sp) begin
                  mem_7 <= io_din;
                end
              end
            end else begin
              mem_7 <= mem_6;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h7 == wr_sp) begin
              mem_7 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_8 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h8 == wr_sp) begin
            mem_8 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_8 <= mem_7;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h8 == wr_sp) begin
                      mem_8 <= io_din;
                    end
                  end
                end else begin
                  mem_8 <= mem_7;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h8 == wr_sp) begin
                  mem_8 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_8 <= mem_7;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_8 <= mem_7;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h8 == wr_sp) begin
                  mem_8 <= io_din;
                end
              end
            end else begin
              mem_8 <= mem_7;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h8 == wr_sp) begin
              mem_8 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_9 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'h9 == wr_sp) begin
            mem_9 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_9 <= mem_8;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'h9 == wr_sp) begin
                      mem_9 <= io_din;
                    end
                  end
                end else begin
                  mem_9 <= mem_8;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'h9 == wr_sp) begin
                  mem_9 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_9 <= mem_8;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_9 <= mem_8;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'h9 == wr_sp) begin
                  mem_9 <= io_din;
                end
              end
            end else begin
              mem_9 <= mem_8;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'h9 == wr_sp) begin
              mem_9 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_10 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'ha == wr_sp) begin
            mem_10 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_10 <= mem_9;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'ha == wr_sp) begin
                      mem_10 <= io_din;
                    end
                  end
                end else begin
                  mem_10 <= mem_9;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'ha == wr_sp) begin
                  mem_10 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_10 <= mem_9;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_10 <= mem_9;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'ha == wr_sp) begin
                  mem_10 <= io_din;
                end
              end
            end else begin
              mem_10 <= mem_9;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'ha == wr_sp) begin
              mem_10 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_11 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'hb == wr_sp) begin
            mem_11 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_11 <= mem_10;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'hb == wr_sp) begin
                      mem_11 <= io_din;
                    end
                  end
                end else begin
                  mem_11 <= mem_10;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'hb == wr_sp) begin
                  mem_11 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_11 <= mem_10;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_11 <= mem_10;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'hb == wr_sp) begin
                  mem_11 <= io_din;
                end
              end
            end else begin
              mem_11 <= mem_10;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'hb == wr_sp) begin
              mem_11 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_12 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'hc == wr_sp) begin
            mem_12 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_12 <= mem_11;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'hc == wr_sp) begin
                      mem_12 <= io_din;
                    end
                  end
                end else begin
                  mem_12 <= mem_11;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'hc == wr_sp) begin
                  mem_12 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_12 <= mem_11;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_12 <= mem_11;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'hc == wr_sp) begin
                  mem_12 <= io_din;
                end
              end
            end else begin
              mem_12 <= mem_11;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'hc == wr_sp) begin
              mem_12 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_13 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'hd == wr_sp) begin
            mem_13 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_13 <= mem_12;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'hd == wr_sp) begin
                      mem_13 <= io_din;
                    end
                  end
                end else begin
                  mem_13 <= mem_12;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'hd == wr_sp) begin
                  mem_13 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_13 <= mem_12;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_13 <= mem_12;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'hd == wr_sp) begin
                  mem_13 <= io_din;
                end
              end
            end else begin
              mem_13 <= mem_12;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'hd == wr_sp) begin
              mem_13 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_14 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'he == wr_sp) begin
            mem_14 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_14 <= mem_13;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'he == wr_sp) begin
                      mem_14 <= io_din;
                    end
                  end
                end else begin
                  mem_14 <= mem_13;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'he == wr_sp) begin
                  mem_14 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_14 <= mem_13;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_14 <= mem_13;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'he == wr_sp) begin
                  mem_14 <= io_din;
                end
              end
            end else begin
              mem_14 <= mem_13;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'he == wr_sp) begin
              mem_14 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      mem_15 <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          if (4'hf == wr_sp) begin
            mem_15 <= io_din;
          end else begin
            if (_T_6) begin
              if (_T_7) begin
                mem_15 <= mem_14;
              end else begin
                if (_T_10) begin
                  if (_T_2) begin
                    if (4'hf == wr_sp) begin
                      mem_15 <= io_din;
                    end
                  end
                end else begin
                  mem_15 <= mem_14;
                end
              end
            end else begin
              if (_T_2) begin
                if (4'hf == wr_sp) begin
                  mem_15 <= io_din;
                end
              end
            end
          end
        end else begin
          mem_15 <= mem_14;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            mem_15 <= mem_14;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                if (4'hf == wr_sp) begin
                  mem_15 <= io_din;
                end
              end
            end else begin
              mem_15 <= mem_14;
            end
          end
        end else begin
          if (_T_2) begin
            if (4'hf == wr_sp) begin
              mem_15 <= io_din;
            end
          end
        end
      end
    end
    if (reset) begin
      dout_reg <= 8'h0;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          dout_reg <= 8'h0;
        end else begin
          dout_reg <= mem_15;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            dout_reg <= mem_15;
          end else begin
            if (!(_T_10)) begin
              dout_reg <= mem_15;
            end
          end
        end
      end
    end
    empty_reg <= reset | _GEN_174;
    if (reset) begin
      wr_sp <= 4'hf;
    end else begin
      if (_T_13) begin
        if (_T_14) begin
          wr_sp <= _T_4;
        end
      end else begin
        if (_T_6) begin
          if (_T_7) begin
            wr_sp <= _T_9;
          end else begin
            if (_T_10) begin
              if (_T_2) begin
                wr_sp <= _T_4;
              end
            end else begin
              wr_sp <= _T_9;
            end
          end
        end else begin
          if (_T_2) begin
            wr_sp <= _T_4;
          end
        end
      end
    end
  end
endmodule
